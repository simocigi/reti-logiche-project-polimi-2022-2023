-- TB EXAMPLE PFRL 2022-2023

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 35; -- 5 + 3 + 20 + 7   (RST) + (CH2-MEM[1]) + 20 CYCLES + (CH1-MEM[6])
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & "000" & "00000000000000000000" & "0000000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & "111" & "00000000000000000000" & "1111100";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & "101" & "00000000000000000000" & "0111000";
    -- Channel 2 -> MEM[1] -> 162
    -- Channel 1 -> MEM[2] -> 75

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  0 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
                                1 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
                                2 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
                                3 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
                                4 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
                                5 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
                                6 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
                                7 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
                                15 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
                                OTHERS => "00110011"-- (OTHERS => '0')
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
                ASSERT (mem_we = '1' OR mem_we = '0') REPORT "o_mem_we in an unexpected state" SEVERITY failure;
            END IF;
            ASSERT (enable_wire = '1' OR enable_wire = '0') REPORT "o_mem_en in an unexpected state" SEVERITY failure;
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        -- wait for 10000 ns;
        tb_rst <= '1';
        wait until falling_edge(tb_clk);
        tb_rst <= '0';
        wait until falling_edge(tb_clk);
        tb_start <= '1';
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        tb_w <= '0';
        wait until falling_edge(tb_clk);
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        tb_start <= '1';
        tb_w <= '1';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        tb_start <= '0';
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        wait until falling_edge(tb_clk);
        
        ASSERT false REPORT "Simulation Ended! TEST PASSATO (EXAMPLE)" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;
